LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY TB_quicksort_tb IS
END TB_quicksort_tb;

ARCHITECTURE TB_quicksort_tb_RTL OF TB_quicksort_tb IS

SIGNAL sim_okay : BOOLEAN := TRUE;

SIGNAL         AP_CE : STD_LOGIC;
SIGNAL        AP_CLK : STD_LOGIC;
SIGNAL        AP_RST : STD_LOGIC;
SIGNAL       DATA_Q0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL        LEFT_R : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL       RIGHT_R : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL DATA_ADDRESS0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL      DATA_CE0 : STD_LOGIC;
SIGNAL       DATA_D0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL      DATA_WE0 : STD_LOGIC;
SIGNAL   OP_PROPERTY : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL  OP_TIMEPOINT : STD_LOGIC_VECTOR(1 DOWNTO 0);

COMPONENT QUICKSORT PORT(
	        AP_CE : IN STD_LOGIC;
	       AP_CLK : IN STD_LOGIC;
	       AP_RST : IN STD_LOGIC;
	      DATA_Q0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	       LEFT_R : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	      RIGHT_R : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DATA_ADDRESS0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
	     DATA_CE0 : OUT STD_LOGIC;
	      DATA_D0 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	     DATA_WE0 : OUT STD_LOGIC;
	  OP_PROPERTY : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	 OP_TIMEPOINT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	 );
END COMPONENT;

BEGIN

DO_SIMULATE: PROCESS
BEGIN

WAIT FOR 0 ns;

	       ap_clk <= '1';
	        ap_ce <= '1';
	       ap_rst <= '1';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 5 ns; 
	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '1';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "10011001000101111111111111111110";
	      right_r <= "10011001000101111111111111111111";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "10011001000101111111111111111110";
	      right_r <= "10011001000101111111111111111111";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00001011001100001000000011000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00001011001100001000000011000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00001011001100001000000011000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00001011001100001000000011000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00001011001100001000000011000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00001011001100001000000011000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11100000110000001000000010100001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010100000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010100000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11000000010100000010110110100000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11000000010100000010110110100000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11000000010100000010110110100000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "11000000010100000010110110100000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100011010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100011010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100011010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100011010111100010110011100101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100110001000010100101100001100";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100110001000010100101100001100";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100100000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100100000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01101000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01101000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100110001000010100101100001100";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100110001000010100101100001100";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100110001000010100101100001100";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100110001000010100101100001100";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100010001000010100101100001101";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100011000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100011000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01101000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01101000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100111010000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100111010000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100111100000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100111100000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01110000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "01011111101011000101010111111111";
	      right_r <= "01011111101011000101011000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "01011111101011000101010111111111";
	      right_r <= "01011111101011000101011000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01011010110011111011110011110001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01011010110011111011110011110001";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01011010110011111100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01011010110011111100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01111100000000000100000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "10000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "01100000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '0';

WAIT FOR 1 ns;

	        ap_ce <= '1';
	       ap_rst <= '0';
	      data_q0 <= "00000000000000000000000000000000";
	       left_r <= "00000000000000000000000000000000";
	      right_r <= "00000000000000000000000000000000";

WAIT FOR 4 ns; 



	       ap_clk <= '1';



END PROCESS;

DUT : QUICKSORT PORT MAP(
	        AP_CE=>AP_CE,
	       AP_CLK=>AP_CLK,
	       AP_RST=>AP_RST,
	      DATA_Q0=>DATA_Q0,
	       LEFT_R=>LEFT_R,
	      RIGHT_R=>RIGHT_R,
	DATA_ADDRESS0=>DATA_ADDRESS0,
	     DATA_CE0=>DATA_CE0,
	      DATA_D0=>DATA_D0,
	     DATA_WE0=>DATA_WE0
	       ,

	     
	  OP_PROPERTY=>OP_PROPERTY,
	 OP_TIMEPOINT=>OP_TIMEPOINT
	 );

END TB_quicksort_tb_RTL;
